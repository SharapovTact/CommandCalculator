library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity const_MODC_Display is
    Port ( MODC : out  STD_LOGIC_VECTOR (9 downto 0));
end const_MODC_Display;

architecture Behavioral of const_MODC_Display is

begin
	MODC <= "1010000000";
end Behavioral;

