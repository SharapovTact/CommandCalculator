library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity const_MODC_PulseWidth is
    Port ( MODC : out  STD_LOGIC_VECTOR (9 downto 0));
end const_MODC_PulseWidth;

architecture Behavioral of const_MODC_PulseWidth is

begin
	MODC <= "0001100000";
end Behavioral;

